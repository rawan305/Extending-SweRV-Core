// NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE
// This is an automatically generated file by nimrodb on Sat Sep 19 23:08:35 IDT 2020
//
// cmd:    swerv -target=default 
//

`include "common_defines.vh"
`undef ASSERT_ON
`undef TEC_RV_ICG
`define TEC_RV_ICG HDBLVT16_CKGTPLT_V5_12
`define PHYSICAL 1
